LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY WriteBackStage IS
	PORT (
		EX_OUT, MEM_OUT  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RDST_INDEX_IN: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
		WRITEDATA  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RDST_INDEX_OUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        REG_WRITE_ENABLE, PORT_WRITE_ENABLE : OUT STD_LOGIC);
END WriteBackStage;

ARCHITECTURE arch_WriteBackStage OF WriteBackStage IS
BEGIN
	WRITEDATA <= EX_OUT WHEN CTRL_SIG_IN(4) = '0'
    ELSE MEM_OUT;

    REG_WRITE_ENABLE <= CTRL_SIG_IN(3);
    PORT_WRITE_ENABLE <= CTRL_SIG_IN(2);
END arch_WriteBackStage;