
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Main IS
        PORT (
        CLK,Reset : IN STD_LOGIC;
        INPUT_PORT : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        OUTPUT_PORT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
END Main;

ARCHITECTURE arch_main OF Main IS

----------------------
----------------------
-- MAIN SIGNALS
----------------------
----------------------

PC, OUTPUT_PORT : STD_LOGIC_VECTOR(31 DOWNTO 0);



----------------------
----------------------
-- STAGES
----------------------
----------------------

COMPONENT FetchStage IS
        PORT (
        CLK : IN STD_LOGIC;
        PC_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        PC_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        INSTRUCTION : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        IMMEDIATE_VALUE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
        );
END COMPONENT;

COMPONENT ExecutionStage IS
	PORT (
		RST : IN STD_LOGIC;
		RSRC_VAL, RDST_VAL, IN_PORT  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RSRC_SHIFT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
		EX_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END COMPONENT;

COMPONENT DecodeStage IS
    PORT (
    CLK: IN STD_LOGIC;
    INSTRUCTION_IN, IMMEDIATE_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    PC_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

    RSRC_INDEX_OUT, RDST_INDEX_OUT : OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
    IMMEDIATE_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); 
    CTRL_SIG : OUT STD_LOGIC_VECTOR(20 DOWNTO 0);
    PC_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;

COMPONENT MemoryStage IS
        PORT (
        -- INPUTS
        CLK : IN STD_LOGIC;
        PC_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        SP_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        Rsrc_value_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        Rdst_value_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        Rsrc_index_IN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        Rdst_index_IN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        Control_Signals_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        ALU_Output_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        -- OUTPUTS
        PC_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        SP_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        Rdst_index_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        ALU_Output_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        MemOutput_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        Control_Signals_OUT : OUT STD_LOGIC_VECTOR(20 DOWNTO 0)
        );
END COMPONENT;

----------------------
----------------------
-- BUFFERS
----------------------
----------------------

COMPONENT IF_ID IS
	PORT (
		CLK, RST, WRITE_ENABLE : IN STD_LOGIC;
		PC_IN  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        INSTRUCTION_IN, IMMEDIATE_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		PC_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        INSTRUCTION_OUT, IMMEDIATE_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT;

COMPONENT ID_EX IS
	PORT (
		CLK, RST, WRITE_ENABLE : IN STD_LOGIC;
		PC_IN, RSRC_VAL_IN, RDST_VAL_IN  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        RSRC_INDEX_IN, RDST_INDEX_IN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		PC_OUT, RSRC_VAL_OUT, RDST_VAL_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RSRC_INDEX_OUT, RDST_INDEX_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        CTRL_SIG_OUT : OUT STD_LOGIC_VECTOR(20 DOWNTO 0));
END COMPONENT;

COMPONENT EX_MEM IS
	PORT (
		CLK, RST, WRITE_ENABLE : IN STD_LOGIC;
		PC_IN, RSRC_VAL_IN, RDST_VAL_IN, EX_IN  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        RSRC_INDEX_IN, RDST_INDEX_IN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		PC_OUT, RSRC_VAL_OUT, RDST_VAL_OUT, EX_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RSRC_INDEX_OUT, RDST_INDEX_OUT  : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        CTRL_SIG_OUT : OUT STD_LOGIC_VECTOR(20 DOWNTO 0));
END COMPONENT;

COMPONENT MEM_WB IS
	PORT (
		CLK, RST, WRITE_ENABLE : IN STD_LOGIC;
		PC_IN, EX_IN, MEM_IN   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        RDST_INDEX_IN  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		PC_OUT, EX_OUT, MEM_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RDST_INDEX_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        CTRL_SIG_OUT : OUT STD_LOGIC_VECTOR(20 DOWNTO 0));
END COMPONENT;

----------------------
----------------------
-- REGISTER FILES
----------------------
----------------------


COMPONENT RegisterFile IS
	GENERIC (N : INTEGER := 32);
	PORT (
		CLK, RST, ENABLE : IN STD_LOGIC;
		InputBus : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        writeIndex, readIndex1, readIndex2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		OutputBus1, OutputBus2 : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0));
END COMPONENT;

    
BEGIN
    
    -- PORTMAPS
    FetchStage_PORTMAP: FetchStage PORT MAP(
        CLK,
        PC,
        PC_OUT,
        INSTRUCTION,
        IMMEDIATE_VALUE
    );

END arch_main;