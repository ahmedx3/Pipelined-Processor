LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY ExecutionStage IS
	PORT (
		CLK, RST : IN STD_LOGIC;
		RSRC_VAL, RDST_VAL, IN_PORT  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RSRC_SHIFT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        DATA_FORWARD_EN_RSRC, DATA_FORWARD_EN_RDST: IN STD_LOGIC;
		DATA_FORWARD_RSRC, DATA_FORWARD_RDST: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RSRC_VAL_EX, RDST_VAL_EX, EX_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        BRANCH : OUT STD_LOGIC;
        BRANCH_VALUE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END ExecutionStage;

ARCHITECTURE arch_ExecutionStage OF ExecutionStage IS
COMPONENT ALU IS
    GENERIC (n : integer:=32);
    PORT ( CLK : IN STD_LOGIC; 
        A,B: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
        SEL: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        SHIFT: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
        FLAG : INOUT STD_LOGIC_VECTOR (2 DOWNTO 0);
        C : OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0);
        FLAG_EN,RST : IN STD_LOGIC);
END COMPONENT;
    SIGNAL FLAG : STD_LOGIC_VECTOR (2 DOWNTO 0) := "000";
    SIGNAL A,B, ALU_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    CONSTANT ZERO : STD_LOGIC_VECTOR (15 DOWNTO 0):=(OTHERS => '0');
BEGIN
	A <= IN_PORT WHEN CTRL_SIG_IN(14 DOWNTO 13) = "11"
    ELSE ZERO & IMMEDIATE WHEN CTRL_SIG_IN(14 DOWNTO 13) = "01"
    ELSE DATA_FORWARD_RSRC WHEN DATA_FORWARD_EN_RSRC = '1'
    ELSE RSRC_VAL WHEN (CTRL_SIG_IN(14 DOWNTO 13) = "00" OR CTRL_SIG_IN(14 DOWNTO 13) = "10") AND DATA_FORWARD_EN_RSRC = '0';
	
    B <= ZERO & IMMEDIATE WHEN CTRL_SIG_IN(14 DOWNTO 13) = "10"
    ELSE DATA_FORWARD_RDST WHEN DATA_FORWARD_EN_RDST = '1'
    ELSE RDST_VAL WHEN (CTRL_SIG_IN(14 DOWNTO 13) = "00" OR CTRL_SIG_IN(14 DOWNTO 13) = "01" OR CTRL_SIG_IN(14 DOWNTO 13) = "11") AND DATA_FORWARD_EN_RDST = '0';

    RSRC_VAL_EX <= DATA_FORWARD_RSRC WHEN DATA_FORWARD_EN_RSRC = '1'
    ELSE RSRC_VAL;

    RDST_VAL_EX <= DATA_FORWARD_RDST WHEN DATA_FORWARD_EN_RDST = '1'
    ELSE RDST_VAL;

    alu0: ALU GENERIC MAP(32) PORT MAP(CLK, A,B,CTRL_SIG_IN(18 DOWNTO 15), RSRC_SHIFT, FLAG, ALU_OUT, CTRL_SIG_IN(8), RST);

    EX_OUT <= ALU_OUT; --NEEDS MODIFICATIONS 

    BRANCH_VALUE <= DATA_FORWARD_RDST WHEN DATA_FORWARD_EN_RDST = '1'
    ELSE RDST_VAL;

    BRANCH <= '1' WHEN CTRL_SIG_IN(20 DOWNTO 19) = "10" AND ( (FLAG(0) = '1' AND CTRL_SIG_IN(2 DOWNTO 1) = "11") OR (FLAG(1) = '1' AND CTRL_SIG_IN(2 DOWNTO 1) = "01") OR (FLAG(2) = '1' AND CTRL_SIG_IN(2 DOWNTO 1) = "10") OR ( CTRL_SIG_IN(2 DOWNTO 1) = "00")  )
    ELSE '0';
END arch_ExecutionStage;