LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY ExecutionStage IS
	PORT (
		RST : IN STD_LOGIC;
		RSRC_VAL, RDST_VAL, IN_PORT  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RSRC_SHIFT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
		EX_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END ExecutionStage;

ARCHITECTURE arch_ExecutionStage OF ExecutionStage IS
COMPONENT ALU IS
    GENERIC (n : integer:=32);
    PORT ( A,B: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
        SEL: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        SHIFT: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
        FLAG : INOUT STD_LOGIC_VECTOR (2 DOWNTO 0);
        C : OUT STD_LOGIC_VECTOR (n-1 DOWNTO 0);
        FLAG_EN,RST : IN STD_LOGIC);
END COMPONENT;
    SIGNAL FLAG : STD_LOGIC_VECTOR (2 DOWNTO 0) := "000";
    SIGNAL A,B, ALU_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
    CONSTANT ZERO : STD_LOGIC_VECTOR (15 DOWNTO 0):=(OTHERS => '0');
BEGIN
	A <= RSRC_VAL WHEN CTRL_SIG_IN(14 DOWNTO 13) = "00" OR CTRL_SIG_IN(14 DOWNTO 13) = "10"
    ELSE ZERO & IMMEDIATE WHEN CTRL_SIG_IN(14 DOWNTO 13) = "01"
    ELSE IN_PORT WHEN CTRL_SIG_IN(14 DOWNTO 13) = "11";
	
    B <= RDST_VAL WHEN CTRL_SIG_IN(14 DOWNTO 13) = "00" OR CTRL_SIG_IN(14 DOWNTO 13) = "01" OR CTRL_SIG_IN(14 DOWNTO 13) = "11"
    ELSE ZERO & IMMEDIATE WHEN CTRL_SIG_IN(14 DOWNTO 13) = "10";

    alu0: ALU GENERIC MAP(32) PORT MAP(A,B,CTRL_SIG_IN(18 DOWNTO 15), RSRC_SHIFT, FLAG, ALU_OUT, CTRL_SIG_IN(8), RST);

    EX_OUT <= ALU_OUT; --NEEDS MODIFICATIONS 
END arch_ExecutionStage;