LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY mREGISTER IS
	GENERIC (N : INTEGER := 32);
	PORT (
		CLK, RST, ENABLE : IN STD_LOGIC;
		D : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
		Q : OUT STD_LOGIC_VECTOR(N - 1 DOWNTO 0));
END mREGISTER;

ARCHITECTURE arch_register OF mREGISTER IS

BEGIN

	PROCESS (CLK, ENABLE, RST)
	BEGIN
		IF RST = '1' THEN
			Q <= (OTHERS => '0');
		ELSIF rising_edge(CLK) AND ENABLE = '1' THEN
			Q <= D;
		END IF;
	END PROCESS;
END arch_register;