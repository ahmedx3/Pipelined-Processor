LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY MEM_WB IS
	PORT (
		CLK, RST, WRITE_ENABLE : IN STD_LOGIC;
		PC_IN, EX_IN, MEM_IN   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        RDST_INDEX_IN  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		PC_OUT, EX_OUT, MEM_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RDST_INDEX_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        CTRL_SIG_OUT : OUT STD_LOGIC_VECTOR(20 DOWNTO 0));
END MEM_WB;

ARCHITECTURE arch_MEM_WB OF MEM_WB IS
BEGIN
	PROCESS (CLK, WRITE_ENABLE, RST)
	BEGIN
		IF RST = '1' THEN
			PC_OUT          <= (OTHERS => '0');
			EX_OUT          <= (OTHERS => '0');
			MEM_OUT         <= (OTHERS => '0');
            RDST_INDEX_OUT  <= (OTHERS => '0');
			CTRL_SIG_OUT    <= (OTHERS => '0');
		ELSIF rising_edge(CLK) AND WRITE_ENABLE = '1' THEN
			PC_OUT          <= PC_IN;
            EX_OUT          <= EX_IN;
			MEM_OUT         <= MEM_IN;
            RDST_INDEX_OUT  <= RDST_INDEX_IN;
			CTRL_SIG_OUT    <=   CTRL_SIG_IN;
		END IF;
	END PROCESS;
END arch_MEM_WB;