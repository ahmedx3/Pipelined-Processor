LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY DataForward IS
	PORT (
		REG_WRITE_EX, REG_WRITE_MEM, MEM_TO_REG : IN STD_LOGIC;
		RDST_INDEX_EX, RDST_INDEX_MEM, RSRC_INDEX_ID, RDST_INDEX_ID : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		ALU_OUT_EX, ALU_OUT_MEM, MEM_OUT_MEM: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_FORWARD_EN_RSRC, DATA_FORWARD_EN_RDST: OUT STD_LOGIC;
		DATA_FORWARD_OUT_RSRC, DATA_FORWARD_OUT_RDST: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END DataForward;

ARCHITECTURE arch_DataForward OF DataForward IS
BEGIN

DATA_FORWARD_EN_RSRC <= '1' WHEN (REG_WRITE_EX = '1' AND RSRC_INDEX_ID = RDST_INDEX_EX) OR (REG_WRITE_MEM = '1' AND RSRC_INDEX_ID = RDST_INDEX_MEM)
ELSE '0';

DATA_FORWARD_EN_RDST <= '1' WHEN (REG_WRITE_EX = '1' AND RDST_INDEX_ID = RDST_INDEX_EX) OR (REG_WRITE_MEM = '1' AND RDST_INDEX_ID = RDST_INDEX_MEM)
ELSE '0';


DATA_FORWARD_OUT_RSRC <= ALU_OUT_EX WHEN (REG_WRITE_EX = '1' AND RSRC_INDEX_ID = RDST_INDEX_EX)
ELSE ALU_OUT_MEM WHEN (REG_WRITE_MEM = '1' AND RSRC_INDEX_ID = RDST_INDEX_MEM) AND MEM_TO_REG = '0'
ELSE MEM_OUT_MEM WHEN (REG_WRITE_MEM = '1' AND RSRC_INDEX_ID = RDST_INDEX_MEM) AND MEM_TO_REG = '1'
ELSE (OTHERS => '0');

DATA_FORWARD_OUT_RDST <= ALU_OUT_EX WHEN (REG_WRITE_EX = '1' AND RDST_INDEX_ID = RDST_INDEX_EX)
ELSE ALU_OUT_MEM WHEN (REG_WRITE_MEM = '1' AND RDST_INDEX_ID = RDST_INDEX_MEM) AND MEM_TO_REG = '0'
ELSE MEM_OUT_MEM WHEN (REG_WRITE_MEM = '1' AND RDST_INDEX_ID = RDST_INDEX_MEM) AND MEM_TO_REG = '1'
ELSE (OTHERS => '0');

END arch_DataForward;