LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY ID_EX IS
	PORT (
		CLK, RST, WRITE_ENABLE, LOAD_USE_STALL : IN STD_LOGIC;
		PC_IN, RSRC_VAL_IN, RDST_VAL_IN  : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        CTRL_SIG_IN : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
        RSRC_INDEX_IN, RDST_INDEX_IN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		PC_OUT, RSRC_VAL_OUT, RDST_VAL_OUT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RSRC_INDEX_OUT, RDST_INDEX_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        IMMEDIATE_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        CTRL_SIG_OUT : OUT STD_LOGIC_VECTOR(20 DOWNTO 0));
END ID_EX;

ARCHITECTURE arch_ID_EX OF ID_EX IS
BEGIN
	PROCESS (CLK, WRITE_ENABLE, RST)
	BEGIN
		IF RST = '1' OR (LOAD_USE_STALL = '1' AND RISING_EDGE(CLK)) THEN
			PC_OUT <= (OTHERS => '0');
			RSRC_VAL_OUT    <= (OTHERS => '0');
			RDST_VAL_OUT    <= (OTHERS => '0');
            RSRC_INDEX_OUT  <= (OTHERS => '0');
            RDST_INDEX_OUT  <= (OTHERS => '0');
			IMMEDIATE_OUT   <= (OTHERS => '0');
			CTRL_SIG_OUT    <= (OTHERS => '0');
		ELSIF rising_edge(CLK) AND WRITE_ENABLE = '1' THEN
			PC_OUT <= PC_IN;
			RSRC_VAL_OUT    <=   RSRC_VAL_IN;
			RDST_VAL_OUT    <=   RDST_VAL_IN;
            RSRC_INDEX_OUT  <= RSRC_INDEX_IN;
            RDST_INDEX_OUT  <= RDST_INDEX_IN;
			IMMEDIATE_OUT   <=  IMMEDIATE_IN;
			CTRL_SIG_OUT    <=   CTRL_SIG_IN;
		END IF;
	END PROCESS;
END arch_ID_EX;